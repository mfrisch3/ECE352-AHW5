module segBdec
(
	input [3:0] D,
	output segB
);

  //////////////////////////////////////////
  // Declare any needed internal signals //
  ////////////////////////////////////////
  logic n1;
  
  //////////////////////////////////////////////////////
  // Write STRUCTURAL verilog to implement segment B //
  ////////////////////////////////////////////////////
  xor iXOR1(n1,D[0],D[1]);
  and iAND1(segB,n1,D[2]);
  
endmodule
